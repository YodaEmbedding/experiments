module hello_world;

initial begin
    $display ("Hello, world!");
    #10 $finish;
end

endmodule
